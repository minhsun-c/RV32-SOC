`include "defines.v"

module id (
    input rst_i,

    //from if_id
    input [`ADDR_WIDTH-1:0] inst_addr_i,
    input [`DATA_WIDTH-1:0] inst_i,

    //from regfile
    input [`RDATA_WIDTH-1:0] reg1_rdata_i,
    input [`RDATA_WIDTH-1:0] reg2_rdata_i,

    // to regfile
    output reg [`RADDR_WIDTH-1:0] reg1_raddr_o,
    output reg [`RADDR_WIDTH-1:0] reg2_raddr_o,
    output reg                    reg1_re_o,
    output reg                    reg2_re_o,

    //to id_exe
    output reg [ `DATA_WIDTH-1:0] inst_o,
    output reg [`RDATA_WIDTH-1:0] op1_o,
    output reg [`RDATA_WIDTH-1:0] op2_o,
    output reg                    reg_we_o,
    output reg [`RADDR_WIDTH-1:0] reg_waddr_o,

    // from FW unit
    input                    fw_en1_o,
    input                    fw_en2_o,
    input [`RDATA_WIDTH-1:0] fw_data1_o,
    input [`RDATA_WIDTH-1:0] fw_data2_o
);

    reg  [`RDATA_WIDTH-1:0] op1_o_final;
    reg  [`RDATA_WIDTH-1:0] op2_o_final;
    wire [             6:0] funct7 = inst_i[31:25];
    wire [             6:0] opcode = inst_i[6:0];
    wire [             2:0] funct3 = inst_i[14:12];

    wire [             4:0] rd = inst_i[11:7];
    wire [             4:0] rs1 = inst_i[19:15];
    wire [             4:0] rs2 = inst_i[24:20];

    // Type-I decode
    wire [`RADDR_WIDTH-1:0] i_reg1_raddr_o;
    wire [`RADDR_WIDTH-1:0] i_reg2_raddr_o;
    wire                    i_reg1_re_o;
    wire                    i_reg2_re_o;
    wire [`RDATA_WIDTH-1:0] i_op1_o;
    wire [`RDATA_WIDTH-1:0] i_op2_o;
    wire                    i_reg_we_o;
    wire [`RADDR_WIDTH-1:0] i_reg_waddr_o;

    id_type_i inst_type_i (
        .inst_i      (inst_i),
        .reg1_rdata_i(reg1_rdata_i),
        .reg1_raddr_o(i_reg1_raddr_o),
        .reg2_raddr_o(i_reg2_raddr_o),
        .reg1_re_o   (i_reg1_re_o),
        .reg2_re_o   (i_reg2_re_o),
        .op1_o       (i_op1_o),
        .op2_o       (i_op2_o),
        .reg_we_o    (i_reg_we_o),
        .reg_waddr_o (i_reg_waddr_o)
    );

    // Type-R decode
    wire [`RADDR_WIDTH-1:0] r_reg1_raddr_o;
    wire [`RADDR_WIDTH-1:0] r_reg2_raddr_o;
    wire                    r_reg1_re_o;
    wire                    r_reg2_re_o;
    wire [`RDATA_WIDTH-1:0] r_op1_o;
    wire [`RDATA_WIDTH-1:0] r_op2_o;
    wire                    r_reg_we_o;
    wire [`RADDR_WIDTH-1:0] r_reg_waddr_o;
    id_type_r inst_type_r (
        .inst_i      (inst_i),
        .reg1_rdata_i(reg1_rdata_i),
        .reg2_rdata_i(reg2_rdata_i),
        .reg1_raddr_o(r_reg1_raddr_o),
        .reg2_raddr_o(r_reg2_raddr_o),
        .reg1_re_o   (r_reg1_re_o),
        .reg2_re_o   (r_reg2_re_o),
        .op1_o       (r_op1_o),
        .op2_o       (r_op2_o),
        .reg_we_o    (r_reg_we_o),
        .reg_waddr_o (r_reg_waddr_o)
    );

    always @(*) begin
        if (rst_i) begin
            inst_o       = `NOP;
            reg1_raddr_o = `ZERO_REG;
            reg2_raddr_o = `ZERO_REG;
            reg1_re_o    = `READ_DISABLE;
            reg2_re_o    = `READ_DISABLE;
            reg_we_o     = `WRITE_DISABLE;
            reg_waddr_o  = `ZERO_REG;
            op1_o_final  = `ZERO;
            op2_o_final  = `ZERO;
        end else begin
            case (opcode)
                `INST_TYPE_I: begin
                    inst_o       = inst_i;
                    reg1_raddr_o = i_reg1_raddr_o;
                    reg2_raddr_o = i_reg2_raddr_o;
                    reg1_re_o    = i_reg1_re_o;
                    reg2_re_o    = i_reg2_re_o;
                    op1_o_final  = i_op1_o;
                    op2_o_final  = i_op2_o;
                    reg_we_o     = i_reg_we_o;
                    reg_waddr_o  = i_reg_waddr_o;
                end
                `INST_TYPE_R_M: begin
                    inst_o       = inst_i;
                    reg1_raddr_o = r_reg1_raddr_o;
                    reg2_raddr_o = r_reg2_raddr_o;
                    reg1_re_o    = r_reg1_re_o;
                    reg2_re_o    = r_reg2_re_o;
                    op1_o_final  = r_op1_o;
                    op2_o_final  = r_op2_o;
                    reg_we_o     = r_reg_we_o;
                    reg_waddr_o  = r_reg_waddr_o;
                end
                `INST_TYPE_LUI: begin
                    inst_o       = inst_i;
                    reg1_raddr_o = `ZERO_REG;
                    reg2_raddr_o = `ZERO_REG;
                    reg1_re_o    = `READ_DISABLE;
                    reg2_re_o    = `READ_DISABLE;
                    op1_o_final  = {inst_i[31:12], {12{1'b0}}};
                    op2_o_final  = `ZERO;
                    reg_we_o     = `WRITE_ENABLE;
                    reg_waddr_o  = rd;
                end
                `INST_TYPE_AUIPC: begin
                    inst_o       = inst_i;
                    reg1_raddr_o = `ZERO_REG;
                    reg2_raddr_o = `ZERO_REG;
                    reg1_re_o    = `READ_DISABLE;
                    reg2_re_o    = `READ_DISABLE;
                    op1_o_final  = inst_addr_i;
                    op2_o_final  = {inst_i[31:12], {12{1'b0}}};
                    reg_we_o     = `WRITE_ENABLE;
                    reg_waddr_o  = rd;
                end
                `INST_TYPE_S: begin
                    inst_o       = inst_i;
                    reg1_raddr_o = rs1;
                    reg2_raddr_o = rs2;
                    reg1_re_o    = `READ_ENABLE;
                    reg2_re_o    = `READ_ENABLE;
                    op1_o_final  = reg1_rdata_i;
                    op2_o_final  = reg2_rdata_i;
                    reg_we_o     = `WRITE_DISABLE;
                    reg_waddr_o  = `ZERO_REG;
                end
                `INST_TYPE_L: begin
                    inst_o       = inst_i;
                    reg1_raddr_o = rs1;
                    reg2_raddr_o = `ZERO_REG;
                    reg1_re_o    = `READ_ENABLE;
                    reg2_re_o    = `READ_DISABLE;
                    op1_o_final  = reg1_rdata_i;
                    op2_o_final  = `ZERO;
                    reg_we_o     = `WRITE_ENABLE;
                    reg_waddr_o  = rd;
                end
                default: begin
                    inst_o       = `NOP;
                    reg1_raddr_o = `ZERO_REG;
                    reg2_raddr_o = `ZERO_REG;
                    reg1_re_o    = `READ_DISABLE;
                    reg2_re_o    = `READ_DISABLE;
                    reg_we_o     = `WRITE_DISABLE;
                    reg_waddr_o  = `ZERO_REG;
                    op1_o_final  = `ZERO;
                    op2_o_final  = `ZERO;
                end
            endcase
        end
    end

    //determine op1_o
    always @(*) begin
        if (fw_en1_o) begin
            op1_o = fw_data1_o;
        end else begin
            op1_o = op1_o_final;
        end
    end

    //determine op2_o
    always @(*) begin
        if (fw_en2_o) begin
            op2_o = fw_data2_o;
        end else begin
            op2_o = op2_o_final;
        end
    end
endmodule

